library verilog;
use verilog.vl_types.all;
entity Deco_vlg_vec_tst is
end Deco_vlg_vec_tst;
